/*
*   Copyright 2016 Purdue University
*   
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*   
*       http://www.apache.org/licenses/LICENSE-2.0
*   
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by Spike 
*/

`define TRACE_FILE_NAME "trace.log"

import rv32i_types_pkg::*;
module cpu_tracker(
  input logic CLK, wb_stall,
  input word_t instr, pc,
  input opcode_t opcode,
  input logic [2:0] funct3
);
  parameter CPUID = 0;

  integer fptr;
  string instr_mnemonic, output_str;
  logic [2:0] branch_funct, load_funct, store_funct;
  logic [2:0] imm_funct, regreg_funct, system_funct;
  logic [63:0] pc64;
  assign pc64 = {{32{1'b0}}, pc};
  initial begin: INIT_FILE
    fptr = $fopen(`TRACE_FILE_NAME, "w");
  end

  always_comb begin
    case (opcode)
      LUI:          instr_mnemonic = "lui";
      AUIPC:        instr_mnemonic = "auipc";
      JAL:          instr_mnemonic = "jal";
      JALR:         instr_mnemonic = "jalr";
      BRANCH: begin
        case(branch_t'(funct3))
          BEQ:      instr_mnemonic = "beq";
          BNE:      instr_mnemonic = "bne";
          BLT:      instr_mnemonic = "blt";
          BGE:      instr_mnemonic = "bge";
          BLTU:     instr_mnemonic = "bltu";
          BGEU:     instr_mnemonic = "bgeu";
          default:  instr_mnemonic = "xxx";
        endcase
      end
      LOAD: begin
        case(load_t'(funct3))
          LB:       instr_mnemonic = "lb";
          LH:       instr_mnemonic = "lh";
          LW:       instr_mnemonic = "lw";
          LBU:      instr_mnemonic = "lbu";
          LHU:      instr_mnemonic = "lhu";
          default:  instr_mnemonic = "xxx";
        endcase
      end
      STORE: begin
        case(store_t'(funct3))
          SB:       instr_mnemonic = "sb";
          SH:       instr_mnemonic = "sh";
          SW:       instr_mnemonic = "sw";
          default:  instr_mnemonic = "xxx";
        endcase
      end
      IMMED: begin
        case(imm_t'(funct3))
          ADDI:     instr_mnemonic = "addi";
          SLTI:     instr_mnemonic = "slti";
          SLTIU:    instr_mnemonic = "sltiu";
          XORI:     instr_mnemonic = "xori";
          ORI:      instr_mnemonic = "ori";
          ANDI:     instr_mnemonic = "andi";
          SLLI:     instr_mnemonic = "slli";
          SRI: begin
            if (instr[30])
                    instr_mnemonic = "srai";
            else
                    instr_mnemonic = "srli";
          end
          default:  instr_mnemonic = "xxx";
        endcase
      end
      REGREG: begin
        case(regreg_t'(funct3))
          ADDSUB: begin
            if (instr[30])
                    instr_mnemonic = "sub";
            else
                    instr_mnemonic = "add";
          end
          SLL:      instr_mnemonic = "sll";
          SLT:      instr_mnemonic = "slt";
          SLTU:     instr_mnemonic = "sltu";
          XOR:      instr_mnemonic = "xor";
          SR: begin
            if (instr[30])
                    instr_mnemonic = "sra";
            else
                    instr_mnemonic = "srl";
          end
          OR:       instr_mnemonic = "or";
          AND:      instr_mnemonic = "and";
          default:  instr_mnemonic = "xxx";
        endcase
      end
      SYSTEM: begin
        case(system_t'(funct3))
          CSRRW:    instr_mnemonic = "csrrw";
          CSRRS:    instr_mnemonic = "csrrs";
          CSRRC:    instr_mnemonic = "csrrc";
          CSRRWI:   instr_mnemonic = "csrrwi";
          CSRRSI:   instr_mnemonic = "csrrsi";
          CSRRCI:   instr_mnemonic = "csrrci";
          default:  instr_mnemonic = "xxx";
        endcase
      end
      default:  instr_mnemonic = "xxx";
    endcase
  end

  always_ff @ (posedge CLK) begin
    if (!wb_stall && instr != 0) begin
      $sformat(output_str, "core%d: 0x%h (0x%h) %s\n", CPUID, pc64, instr, instr_mnemonic);
      $fwrite(fptr, output_str);
    end
  end

  final begin: CLOSE_FILE
    $fclose(fptr);
  end

endmodule
