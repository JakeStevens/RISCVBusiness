
`include "pipe5_hazard_forwarding_unit_if.vh"
`include "prv_pipeline_if.vh"


module pipe5_hazard_forwarding_unit(
    pipe5_hazard_forwarding_unit_if.hazard_unit hazard_if,
    prv_pipeline_if.hazard prv_pipeline_if
);





endmodule
