/*
*   Copyright 2016 Purdue University
*   
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*   
*       http://www.apache.org/licenses/LICENSE-2.0
*   
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*   
*   
*   Filename:     icache.sv
*   
*   Created by:   John Skubic
*   Email:        jskubic@purdue.edu
*   Date Created: 06/01/2016
*   Description:  Instruction Cache	
*/

`include "ram_if.vh"

module icache (
  input logic CLK, nRST,
  ram_if.cpu mem_ram_if,
  ram_if.ram proc_ram_if
);

  //passthrough layer
  assign mem_ram_if.addr     = proc_ram_if.addr;
  assign mem_ram_if.ren      = proc_ram_if.ren;
  assign mem_ram_if.wen      = proc_ram_if.wen;
  assign mem_ram_if.wdata    = proc_ram_if.wdata;
  assign mem_ram_if.byte_en  = proc_ram_if.byte_en; 

  assign proc_ram_if.rdata   = mem_ram_if.rdata;
  assign proc_ram_if.busy    = mem_ram_if.busy;

endmodule
