package pipe5_types_pkg;

endpackage
