`ifndef TSPP_TYPES_PKG_VH
`define TSPP_TYPES_PKG_VH

// include the packages needed for TSPP
`include "rv32i_types_pkg"

package tspp_types_pkg;
  // import those packages
  import rv32i_types_pkg::*;
endpackage
`endif
