package pipe5_types_pkg;

    typedef enum logic[1:0] {
        NO_FWD,
        FWD_M,
        FWD_W
    } bypass_t;

endpackage
