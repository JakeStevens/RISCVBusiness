
module pipe5();


endmodule
