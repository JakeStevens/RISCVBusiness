/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by Spike
*/

`define TRACE_FILE_NAME "trace.log"

module cpu_tracker (
    input logic CLK, wb_stall, instr_30,
    input rv32i_types_pkg::word_t instr, pc,
    input rv32i_types_pkg::opcode_t opcode,
    input logic [2:0] funct3,
    input logic [11:0] funct12,
    input logic [4:0] rs1, rs2, rd,
    input logic [12:0] imm_SB,
    input logic [11:0] imm_S, imm_I,
    input logic [20:0] imm_UJ,
    input logic [31:0] imm_U
);
    import rv32i_types_pkg::*;
    import machine_mode_types_1_12_pkg::*;

    parameter int CPUID = 0;

    integer fptr;
    string instr_mnemonic, output_str, src1, src2, dest, operands;
    string csr, temp_str;
    logic [63:0] pc64;
    assign pc64 = {{32{1'b0}}, pc};
    initial begin : INIT_FILE
        fptr = $fopen(`TRACE_FILE_NAME, "w");
    end

    always_comb begin
        src1 = registerAssign(rs1);
        src2 = registerAssign(rs2);
        dest = registerAssign(rd);
        csr  = csrRegisterAssign(funct12);
    end

    always_comb begin
        case (opcode)
            LUI, AUIPC: $sformat(operands, "%s, %d", dest, imm_U[31:12]);
            JAL:        $sformat(operands, "%s, pc + %d", dest, signed'(imm_UJ));
            JALR:       $sformat(operands, "%s, %s, %d", dest, src1, signed'(imm_I));
            BRANCH:     $sformat(operands, "%s, %s, pc + %d", src1, src2, signed'(imm_SB));
            STORE:      $sformat(operands, "%s, %d(%s)", src2, signed'(imm_S), src1);
            LOAD:       $sformat(operands, "%s, %d(%s)", dest, signed'(imm_I), src1);
            IMMED:      $sformat(operands, "%s, %s, %d", dest, src1, signed'(imm_I));
            REGREG:     $sformat(operands, "%s, %s, %s", dest, src1, src2);
            SYSTEM: begin
                case (rv32i_system_t'(funct3))
                    CSRRS, CSRRW, CSRRC:    $sformat(operands, "%s, %s, %s", dest, csr, src1);
                    CSRRSI, CSRRWI, CSRRCI: $sformat(operands, "%s, %s, %d", dest, csr, rs1);
                    PRIV:                   operands = "";
                    default:                operands = "";
                endcase
            end
            default:    operands = "";
        endcase
    end

    always_comb begin
        case (opcode)
            LUI:     instr_mnemonic = "lui";
            AUIPC:   instr_mnemonic = "auipc";
            JAL:     instr_mnemonic = "jal";
            JALR:    instr_mnemonic = "jalr";
            BRANCH: begin
                case (branch_t'(funct3))
                    BEQ:     instr_mnemonic = "beq";
                    BNE:     instr_mnemonic = "bne";
                    BLT:     instr_mnemonic = "blt";
                    BGE:     instr_mnemonic = "bge";
                    BLTU:    instr_mnemonic = "bltu";
                    BGEU:    instr_mnemonic = "bgeu";
                    default: instr_mnemonic = "unknown branch op";
                endcase
            end
            LOAD: begin
                case (load_t'(funct3))
                    LB:      instr_mnemonic = "lb";
                    LH:      instr_mnemonic = "lh";
                    LW:      instr_mnemonic = "lw";
                    LBU:     instr_mnemonic = "lbu";
                    LHU:     instr_mnemonic = "lhu";
                    default: instr_mnemonic = "unknown load op";
                endcase
            end
            STORE: begin
                case (store_t'(funct3))
                    SB:      instr_mnemonic = "sb";
                    SH:      instr_mnemonic = "sh";
                    SW:      instr_mnemonic = "sw";
                    default: instr_mnemonic = "unknown store op";
                endcase
            end
            IMMED: begin
                case (imm_t'(funct3))
                    ADDI:    instr_mnemonic = "addi";
                    SLTI:    instr_mnemonic = "slti";
                    SLTIU:   instr_mnemonic = "sltiu";
                    XORI:    instr_mnemonic = "xori";
                    ORI:     instr_mnemonic = "ori";
                    ANDI:    instr_mnemonic = "andi";
                    SLLI:    instr_mnemonic = "slli";
                    SRI: begin
                        if (instr_30) instr_mnemonic = "srai";
                        else instr_mnemonic = "srli";
                    end
                    default: instr_mnemonic = "unknown immed op";
                endcase
            end
            REGREG: begin
                case (regreg_t'(funct3))
                    ADDSUB: begin
                        if (instr_30) instr_mnemonic = "sub";
                        else instr_mnemonic = "add";
                    end
                    SLL:     instr_mnemonic = "sll";
                    SLT:     instr_mnemonic = "slt";
                    SLTU:    instr_mnemonic = "sltu";
                    XOR:     instr_mnemonic = "xor";
                    SR: begin
                        if (instr_30) instr_mnemonic = "sra";
                        else instr_mnemonic = "srl";
                    end
                    OR:      instr_mnemonic = "or";
                    AND:     instr_mnemonic = "and";
                    default: instr_mnemonic = "unknown regreg op";
                endcase
            end
            SYSTEM: begin
                case (rv32i_system_t'(funct3))
                    CSRRW:   instr_mnemonic = "csrrw";
                    CSRRS:   instr_mnemonic = "csrrs";
                    CSRRC:   instr_mnemonic = "csrrc";
                    CSRRWI:  instr_mnemonic = "csrrwi";
                    CSRRSI:  instr_mnemonic = "csrrsi";
                    CSRRCI:  instr_mnemonic = "csrrci";
                    PRIV: begin
                        case (priv_insn_t'(funct12))
                            ECALL:  instr_mnemonic = "ecall";
                            EBREAK: instr_mnemonic = "ebreak";
                            MRET:   instr_mnemonic = "mret";
                            default: begin
                                instr_mnemonic = "errr";
                                $display("%b", priv_insn_t'(funct12));
                            end
                        endcase
                    end
                    default: instr_mnemonic = "unknown system op";
                endcase
            end
            MISCMEM: begin
                case (rv32i_miscmem_t'(funct3))
                    FENCE:   instr_mnemonic = "fence";
                    FENCEI:  instr_mnemonic = "fence.i";
                    default: instr_mnemonic = "unknown misc-mem op";
                endcase
            end
            default: instr_mnemonic = "xxx";
        endcase
    end

    function string registerAssign(input logic [4:0] register);
        case (register)
            5'd0:  registerAssign = "zero";
            5'd1:  registerAssign = "ra";
            5'd2:  registerAssign = "sp";
            5'd3:  registerAssign = "gp";
            5'd4:  registerAssign = "tp";
            5'd5:  registerAssign = "t0";
            5'd6:  registerAssign = "t1";
            5'd7:  registerAssign = "t2";
            5'd8:  registerAssign = "s0";
            5'd9:  registerAssign = "s1";
            5'd10: registerAssign = "a0";
            5'd11: registerAssign = "a1";
            5'd12: registerAssign = "a2";
            5'd13: registerAssign = "a3";
            5'd14: registerAssign = "a4";
            5'd15: registerAssign = "a5";
            5'd16: registerAssign = "a6";
            5'd17: registerAssign = "a7";
            5'd18: registerAssign = "s2";
            5'd19: registerAssign = "s3";
            5'd20: registerAssign = "s4";
            5'd21: registerAssign = "s5";
            5'd22: registerAssign = "s6";
            5'd23: registerAssign = "s7";
            5'd24: registerAssign = "s8";
            5'd25: registerAssign = "s9";
            5'd26: registerAssign = "s10";
            5'd27: registerAssign = "s11";
            5'd28: registerAssign = "t3";
            5'd29: registerAssign = "t4";
            5'd30: registerAssign = "t5";
            5'd31: registerAssign = "t6";
            default: registerAssign = "UNKNOWN REGISTER";
        endcase
    endfunction

    function string csrRegisterAssign(input logic [11:0] csr_register);
        case (csr_addr_t'(csr_register))
            MVENDORID_ADDR: csrRegisterAssign = "mvendorid";
            MARCHID_ADDR:   csrRegisterAssign = "marchid";
            MIMPID_ADDR:    csrRegisterAssign = "mimpid";
            MHARTID_ADDR:   csrRegisterAssign = "mhartid";
            MSTATUS_ADDR:   csrRegisterAssign = "mstatus";
            MISA_ADDR:      csrRegisterAssign = "misa";
            MEDELEG_ADDR:   csrRegisterAssign = "medeleg";
            MIDELEG_ADDR:   csrRegisterAssign = "mideleg";
            MTVEC_ADDR:     csrRegisterAssign = "mtvec";
            MIE_ADDR:       csrRegisterAssign = "mie";
            MSCRATCH_ADDR:  csrRegisterAssign = "mscratch";
            MEPC_ADDR:      csrRegisterAssign = "mepc";
            MCAUSE_ADDR:    csrRegisterAssign = "mcause";
            MTVAL_ADDR:     csrRegisterAssign = "mtval";
            MIP_ADDR:       csrRegisterAssign = "mip";
            default:        csrRegisterAssign = "csr register not tracked";
        endcase
    endfunction

    always_ff @(posedge CLK) begin
        if (!wb_stall && instr != 0) begin
            $sformat(temp_str, "core%d: 0x%h (0x%h)", CPUID, pc64, instr);
            $sformat(output_str, "%s %s %s\n", temp_str, instr_mnemonic, operands);
            $fwrite(fptr, output_str);
        end
    end

    final begin : CLOSE_FILE
        $fclose(fptr);
    end

endmodule
