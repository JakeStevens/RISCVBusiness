`include "ram_if.vh"

module RISCVBusiness (
  input logic CLK, nRST,
  ram_if.cpu ramif
);


endmodule
